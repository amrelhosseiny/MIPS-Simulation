module alu_branch (in1,in2,out1);
input [31:0] in1 ,in2;
output [31:0] out1;

   assign out1=in1+in2;
endmodule
      
     
